LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

ENTITY multiplicador IS
GENERIC (N: INTEGER := 4);
--PORT ();
END multiplicador;

ARCHITECTURE estrutura OF multiplicador IS
BEGIN

END estrutura;